** 4-bit ripple counter
.subckt inverter 1 2 3
.model pmod pmos level=54 version=4.7
.model nmod nmos level=54 version=4.7
mp 2 1 3 3 pmod w=100u l=10u
mn 2 1 0 0 nmod w=100u l=10u
.ends
.subckt dff 1 2 7 8
.model pmod pmos level=54 version=4.7
.model nmod nmos level=54 version=4.7
m1 2 1 3 3 nmod w=100u l=10u
m2 5 1 3 3 pmod w=100u l=10u
m3 6 1 5 5 pmod w=100u l=10u
m4 6 1 8 8 nmod w=100u l=10u
m5 4 3 9 9 pmod w=100u l=10u
m6 4 3 0 0 nmod w=100u l=10u
m7 5 4 9 9 pmod w=100u l=10u
m8 5 4 0 0 nmod w=100u l=10u
m9 7 6 9 9 pmod w=100u l=10u
m10 7 6 0 0 nmod w=100u l=10u
m11 8 7 9 9 pmod w=100u l=10u
m12 8 7 0 0 nmod w=100u l=10u
.ends
Vd 1 0 dc 5v
Vp 11 0 pulse(0 5 0 0 0 10m 20m)
xd1 11 12 12 13 dff
xd2 12 14 14 15 dff
xd3 14 16 16 17 dff
xd4 16 18 18 19 dff
.tran 0.01ms 100ms
.control
run
plot V(11)
plot V(13)
plot V(15)
plot V(17)
plot V(19)
.endc 
.end
